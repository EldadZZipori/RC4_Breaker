`default_nettype none
/*
	KSA
*/

module ksa
(
	input logic CLOCK_50

);
	


endmodule 