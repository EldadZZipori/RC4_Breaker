`default_nettype none
/*
	DECRYPTOR FSM
	This module implements the third loop in the decryption algorithem.
	
	NOTE: This module does not write into S memory! It is ment to be used with a local
			register that is a copy of S memory.
	
	i=0 j = 0
	for k = 0 to key_length-1
		i = i + 1
		j = (j + s[i])
		swap value of s[i] and s[j]
		f = s[ s[i] + s[j]]
		decrypted_output[k] = f xor encrypted_input[k]
		
	This module has three paramters -
	MSG_DEP					number of words in the encrypted data 
	S_DEP						number of words in S memory to be used to crack encryption
	MSG_WIDTH				number of bits in each word (has to be the same in both)
*/

module decryptor_fsm
# (
	parameter MSG_DEP		= 32, 
	parameter S_DEP	 	= 256, 
	parameter MSG_WIDTH 	= 8
)
(
	input logic							clk,
	input logic							reset,
	input logic [MSG_WIDTH-1:0]	encrypted_input[MSG_DEP-1:0],			// the ROM memory containing the encrpted data
	input logic [MSG_WIDTH-1:0]	s_data[S_DEP-1:0],						// locally registred S memory
	input logic [MSG_WIDTH-1:0]	s_q_data_in,
	input logic							start,										// flag indicating this FSM can start operation, Master should insure all other FSM's are done
	
	output logic [MSG_WIDTH-1:0]	address_out,								// Address of local registred S memory to be written to
	output logic [MSG_WIDTH-1:0]	data_out,									// Data to be written to local registred S memory
	output logic 						enable_write,								// Write enable to local registres S memory
	output logic [MSG_WIDTH-1:0]	decrypted_output[MSG_DEP-1:0],		// Decrypted message, to be determined if correct by another FSM
	output logic						done											// Indicates FSM is done operation
);

	/*
		STATE CONTROL
	*/
	localparam IDLE 					= 4'b0000;
	localparam INCREMENT_INDEX_I	= 4'b0011;									// i = i + 1
	localparam INCREMENT_INDEX_J	= 4'b0100;									// j = (j + s[i])
	localparam TAKE_TEMP				= 4'b1111;									// temp = s[j]
	localparam I_TO_J					= 4'b0111;
	localparam WAIT_I_TO_J			= 4'b1001;									// s[j] = s[i]
	localparam DIS_I_TO_J			= 4'b1011;									// This start lowers the enable flag to ensure we are not writing to the wrong address
	localparam J_TO_I					= 4'b1000;
	localparam WAIT_J_TO_I			= 4'b1010;									// s[i] = s[j]
	localparam DIS_J_TO_I			= 4'b1100;									// This start lowers the enable flag to ensure we are not writing to the wrong address
	localparam ASSIGN_F				= 4'b0001;									// f = s[ s[i] + s[j]]
	localparam DECRYPT				= 4'b0010;									// decrypted_output[k] = f xor encrypted_input[k]
	localparam DETERMINE				= 4'b0101;									// k == 255 ? DONE : INCREMENT_INDEX_I
	localparam DONE					= 4'b0110;
	
	
	logic [4:0] current_state/*synthesis keep*/;
	logic [4:0] next_state;
	
	logic [MSG_WIDTH-1:0] 	f;	
	logic	[7:0]					index_i, index_j;
	
	logic [MSG_WIDTH:0] temp_j;
	
	// Flip flop to register the current state
	always_ff @(posedge clk) begin
		current_state <= next_state;
	end
	
	always_comb begin
		if(reset) next_state <= IDLE;
		else begin
			case (current_state)
				IDLE: begin
					if (start) 	next_state <= INCREMENT_INDEX_I;					// Only get out of IDLE start when Master confirmed all other FSM are done execution
					else 			next_state <= IDLE;
					
				end
				INCREMENT_INDEX_I: begin
					next_state = INCREMENT_INDEX_J;
				end
				INCREMENT_INDEX_J: begin
					next_state = TAKE_TEMP;
				end
				TAKE_TEMP: begin
					next_state = I_TO_J;
				end
				I_TO_J: begin
					next_state = WAIT_I_TO_J;
				end
				WAIT_I_TO_J: begin
					next_state = DIS_I_TO_J;
				end
				DIS_I_TO_J: begin
					next_state = J_TO_I;
				end
				J_TO_I: begin
					next_state = WAIT_J_TO_I;
				end
				WAIT_J_TO_I: begin
					next_state = DIS_J_TO_I;
				end
				DIS_J_TO_I: begin
					next_state = ASSIGN_F;
				end
				ASSIGN_F: begin
					next_state = DECRYPT;
				end
				DECRYPT: begin
					next_state = DETERMINE;
				end
				DETERMINE: begin
					if (index_i == ({MSG_WIDTH{1'b1}}))  	next_state = DONE;					// when all data is read stop decryption prosses
					else												next_state = INCREMENT_INDEX_I;	
				end
				DONE: begin
					next_state = DONE;
				end
				default: next_state = IDLE;
			endcase
		end
	end
		
	always_ff @ (posedge clk) begin
		case (current_state)
			IDLE: begin
				index_i 			<= 0;																									
				index_j			<= 0;
				enable_write 	<= 1'b0;
				done 				<= 1'b0;
			end
			INCREMENT_INDEX_I: begin
				index_i <= index_i + 1;
			end
			INCREMENT_INDEX_J: begin
				index_j <= index_j + s_data[index_i];
			end
			TAKE_TEMP: begin
				temp_j <= s_data[index_j];
			end
			I_TO_J: begin
				address_out 	<= index_j;
				data_out			<= s_data[index_i];
				enable_write 	<= 1'b0;
			end
			WAIT_I_TO_J: begin	
				enable_write 	<= 1'b1;
			end
			DIS_I_TO_J: begin
				enable_write 	<= 1'b0;
			end
			J_TO_I: begin
				enable_write 	<= 1'b0;
				address_out 	<= index_i;
				data_out			<= temp_j;
			end
			WAIT_J_TO_I: begin
				enable_write 	<= 1'b1;
			end
			DIS_J_TO_I: begin
				enable_write 	<= 1'b0;
			end
			ASSIGN_F: begin
				f <= s_data[s_data[index_i] +s_data[index_j]];
			end
			DECRYPT: begin
				decrypted_output[index_i-1] <= f ^ encrypted_input[index_i-1]; // k = i -1 always
			end
			DONE: begin
				done <= 1'b1;
			end

		endcase
	end
	
endmodule
